library verilog;
use verilog.vl_types.all;
entity TestBenchProcessor is
end TestBenchProcessor;
