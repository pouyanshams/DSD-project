library verilog;
use verilog.vl_types.all;
entity STACK_BASED_ALU_testbench is
end STACK_BASED_ALU_testbench;
